// See LICENSE.vyoma for more details

module adder(a, b, sum);

 
